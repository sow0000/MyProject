////////////////////////////////////////////////////////////////
//	TITLE : Program Counter
//	FILE : PC.v	
//	ORGANIZATION : Kwangwoon Univ. Computer Engineering
//	STUDENT ID : 2010720092, 2010720117
//	STUDENT NAME : Hyunjae Lee, Seongjoong Kim		
//	PLATFORM : Windows 7
//	SIMULATOR : ModelSim PE Student Edition 10.3	
//	COMPILER : ModelSim PE Student Edition 10.3	
//	DESCRIPTION : This module defines Program Counter.	
//								Use 32 bit Register, and Reset signal.
//	LAST UPDATE : 04.07, 2014
////////////////////////////////////////////////////////////////
module PC(i_next_pc,o_pc,i_rst_n,i_clk,PC_Write);
	input [31:0] i_next_pc;
 	input i_rst_n,i_clk,PC_Write;
	output reg [31:0] o_pc;

	always @ (posedge i_clk or negedge i_rst_n) // clock is rising edge or reset is falling edge
	begin
		if(i_rst_n==0) o_pc <= 32'h0000_0000; // if Reset is ON, then output is 0
		else if(PC_Write==1) o_pc <= i_next_pc; // if Reset is OFF, then output is next pc
		else o_pc <= o_pc;
	end

endmodule
