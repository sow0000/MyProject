////////////////////////////////////////////////////////////////
//	TITLE : 5to32 Decoder
//	FILE : RF_dec532.v	
//	ORGANIZATION : Kwangwoon Univ. Computer Engineering	
//	STUDENT ID : 2010720092, 2010720117	
//	STUDENT NAME : Hyunjae Lee, Seongjoong Kim	
//	PLATFORM : Windows 7	
//	SIMULATOR : ModelSim PE Student Edition 10.3	
//	COMPILER : ModelSim PE Student Edition 10.3	
//	DESCRIPTION : This module defines 5 to 32 Decoder.	
//								Use case function, output each value.
//	LAST UPDATE : 04.07, 2014	
////////////////////////////////////////////////////////////////
module dec532(a,y);
	input [4:0] a;
	output reg [32:0] y;
	
	// Use case function, insert each 32 bit value
	always@(a)
	begin
	case(a)
		5'b00000 : y <= 32'b00000000_00000000_00000000_00000001;
		5'b00001 : y <= 32'b00000000_00000000_00000000_00000010;
		5'b00010 : y <= 32'b00000000_00000000_00000000_00000100;
		5'b00011 : y <= 32'b00000000_00000000_00000000_00001000;
		5'b00100 : y <= 32'b00000000_00000000_00000000_00010000; 
		5'b00101 : y <= 32'b00000000_00000000_00000000_00100000; 
		5'b00110 : y <= 32'b00000000_00000000_00000000_01000000; 
		5'b00111 : y <= 32'b00000000_00000000_00000000_10000000; 
		5'b01000 : y <= 32'b00000000_00000000_00000001_00000000; 
		5'b01001 : y <= 32'b00000000_00000000_00000010_00000000; 
		5'b01010 : y <= 32'b00000000_00000000_00000100_00000000; 
		5'b01011 : y <= 32'b00000000_00000000_00001000_00000000; 
		5'b01100 : y <= 32'b00000000_00000000_00010000_00000000; 
		5'b01101 : y <= 32'b00000000_00000000_00100000_00000000;
		5'b01110 : y <= 32'b00000000_00000000_01000000_00000000;
		5'b01111 : y <= 32'b00000000_00000000_10000000_00000000;
		5'b10000 : y <= 32'b00000000_00000001_00000000_00000000;
		5'b10001 : y <= 32'b00000000_00000010_00000000_00000000;
		5'b10010 : y <= 32'b00000000_00000100_00000000_00000000;
		5'b10011 : y <= 32'b00000000_00001000_00000000_00000000;
		5'b10100 : y <= 32'b00000000_00010000_00000000_00000000;
		5'b10101 : y <= 32'b00000000_00100000_00000000_00000000;
		5'b10110 : y <= 32'b00000000_01000000_00000000_00000000;
		5'b10111 : y <= 32'b00000000_10000000_00000000_00000000;
		5'b11000 : y <= 32'b00000001_00000000_00000000_00000000;
		5'b11001 : y <= 32'b00000010_00000000_00000000_00000000;
		5'b11010 : y <= 32'b00000100_00000000_00000000_00000000;
		5'b11011 : y <= 32'b00001000_00000000_00000000_00000000;
		5'b11100 : y <= 32'b00010000_00000000_00000000_00000000;
		5'b11101 : y <= 32'b00100000_00000000_00000000_00000000;
		5'b11110 : y <= 32'b01000000_00000000_00000000_00000000;
		5'b11111 : y <= 32'b10000000_00000000_00000000_00000000;
	endcase
	end
	
endmodule
